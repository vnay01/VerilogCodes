/*
    Date: 09-feb-2025 :: Vinay Singh
    Testbench for verifying matrix multiplier
*/



