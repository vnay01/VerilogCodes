// N-bit binary Ripple Counter
module udp_ripple_counter(
							output [N-1:0] count_out,
							input count_in, 
							);